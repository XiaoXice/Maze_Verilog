`define MEMORYSIZE 2

module Maze(
  
);

endmodule // MAZE