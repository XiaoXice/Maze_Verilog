module MAZE(
  
);

endmodule // MAZE