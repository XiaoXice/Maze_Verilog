module nvidia(
  input clk; //50MHz
  input [`MEMORYSIZE-1:0] data;
  input []
);

endmodule // nvidia