module commend(
  input clk,
  input key_value,
  output [5:0]address,
  output commend,
  inout [`MEMORYSIZE-1:0] data
);



endmodule // commend