module Maze(
  input clk,
  input nst,
  input [3:0] key_row,
  input [3:0] key_col,
  output [7:0] led_row,
  output [7:0] led_r_col,
  output [7:0] led_g_col
);

endmodule // Maze